/home/013829283/224hw31/EE224_Project/adder1bit/netlist